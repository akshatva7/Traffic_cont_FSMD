
`include "transaction.sv"
`include "generator.sv"
`include "tlc_cov.sv"
`include "tlc_bfm.sv"
`include "intf.sv"

`include "environment.sv"
`include "test.sv"

`include "fsm_d.v"
`include "top.sv"


